module hello_world ;

initial begin
  $display ("Installation successful!");
  #10 $finish;
end

endmodule // End of Module hello_world