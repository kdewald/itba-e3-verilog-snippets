module hello_world ;

initial begin
  $display ("Installation successful!");
  $finish;
end

endmodule // End of Module hello_world